/* verilator lint_off UNUSEDSIGNAL */

module spi_ctrl_top (
    // Clock and resets
    input logic         sys_clk,
    input logic         rst_n
);

endmodule // spi_ctrl_top
