module apb_bridge_tb;

    apb_bridge_top u_apb_bridge_top();

endmodule // apb_bridge_tb
