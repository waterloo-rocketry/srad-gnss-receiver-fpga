module apb_bridge_top;

endmodule // apb_bridge_top
