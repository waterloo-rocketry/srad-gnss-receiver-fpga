/* verilator lint_off PINMISSING */

module periph_subsys_top;

    apb_bridge_top u_apb_bridge_top();

    gpio_ctrl_top u_gpio_ctrl_top();

endmodule // periph_subsys_top
