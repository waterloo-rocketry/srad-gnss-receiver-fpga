module periph_subsys_tb;

    periph_subsys_top u_periph_subsys_top();

endmodule // periph_subsys_tb
